module multipliere();

  reg [7:0]bias1[199:0];
  
  initial begin

	bias1[0]=-40;bias1[1]=-62;bias1[2]=-58;bias1[3]=-12;bias1[4]=-50;bias1[5]=-19;bias1[6]=-52;bias1[7]=-43;bias1[8]=-42;bias1[9]=-71;bias1[10]=-69;bias1[11]=-34;bias1[12]=-26;bias1[13]=-14;bias1[14]=-51;bias1[15]=-28;bias1	[16]=-56;bias1[17]=-47;bias1[18]=-42;bias1[19]=-60;bias1[20]=-40;bias1[21]=-47;bias1[22]=-39;bias1[23]=-67;bias1[24]=-39;bias1[25]=-38;bias1[26]=-48;bias1[27]=-59;bias1[28]=-24;bias1[29]=31;bias1[30]=-22;bias1[31]=-32;bias1[32]=-22;bias1[33]=-34;bias1[34]=-30;bias1[35]=-48;bias1[36]=-19;bias1[37]=-14;bias1[38]=-38;bias1[39]=-42;bias1[40]=-60;bias1[41]=-34;bias1[42]=-67;bias1[43]=-39;bias1[44]=-14;bias1[45]=-45;bias1[46]=-23;bias1[47]=-23;bias1[48]=-28;bias1[49]=-12;bias1[50]=-45;bias1[51]=-17;bias1[52]=-75;bias1[53]=-46;bias1[54]=-63;bias1[55]=-39;bias1[56]=-52;bias1[57]=-73;bias1[58]=-37;bias1[59]=-30;bias1[60]=-16;bias1[61]=-44;bias1[62]=-31;bias1[63]=-73;bias1[64]=-64;bias1[65]=-31;bias1[66]=-59;bias1[67]=-47;bias1[68]=-8;bias1[69]=-20;bias1[70]=-42;bias1[71]=-14;bias1[72]=-73;bias1[73]=-29;bias1[74]=-39;bias1[75]=-47;bias1[76]=-29;bias1[77]=-33;bias1[78]=-31;bias1[79]=-37;bias1[80]=-46;bias1[81]=-65;bias1[82]=-28;bias1[83]=-7;bias1[84]=-52;bias1[85]=-42;bias1[86]=-60;bias1[87]=-33;bias1[88]=-70;bias1[89]=-33;bias1[90]=-36;bias1[91]=-14;bias1[92]=-62;bias1[93]=-34;bias1[94]=-16;bias1[95]=-49;bias1[96]=-36;bias1[97]=-37;bias1[98]=-35;bias1[99]=-49;bias1[100]=-40;bias1[101]=-37;bias1[102]=-54;bias1[103]=-32;bias1[104]=-40;bias1[105]=-23;bias1[106]=-28;bias1[107]=-48;bias1[108]=-28;bias1[109]=-71;bias1[110]=-33;bias1[111]=-34;bias1[112]=-47;bias1[113]=-19;bias1[114]=-21;bias1[115]=-77;bias1[116]=-70;bias1[117]=-14;bias1[118]=-11;bias1[119]=-25;bias1[120]=-31;bias1[121]=-33;bias1[122]=-44;bias1[123]=10;bias1[124]=-21;bias1[125]=-47;bias1[126]=-51;bias1[127]=-57;bias1[128]=-59;bias1[129]=-31;bias1[130]=-28;bias1[131]=-49;bias1[132]=-45;bias1[133]=-10;bias1[134]=-16;bias1[135]=0;bias1[136]=-46;bias1[137]=-31;bias1[138]=-47;bias1[139]=-69;bias1[140]=-41;bias1[141]=-28;bias1[142]=-51;bias1[143]=-14;bias1[144]=-41;bias1[145]=-61;bias1[146]=-52;bias1[147]=-100;bias1[148]=-36;bias1[149]=-27;bias1[150]=-45;bias1[151]=-47;bias1[152]=-19;bias1[153]=-36;bias1[154]=-58;bias1[155]=-85;bias1[156]=-22;bias1[157]=25;bias1[158]=-38;bias1[159]=-61;bias1[160]=-26;bias1[161]=-54;bias1[162]=-27;bias1[163]=-38;bias1[164]=-48;bias1[165]=-42;bias1[166]=-14;bias1[167]=-45;bias1[168]=-19;bias1[169]=-44;bias1[170]=-63;bias1[171]=-22;bias1[172]=-17;bias1[173]=-43;bias1[174]=-33;bias1[175]=-29;bias1[176]=-43;bias1[177]=-71;bias1[178]=-51;bias1[179]=-10;bias1[180]=-49;bias1[181]=-44;bias1[182]=-70;bias1[183]=-39;bias1[184]=-29;bias1[185]=-67;bias1[186]=-38;bias1[187]=-75;bias1[188]=-29;bias1[189]=-61;bias1[190]=-76;bias1[191]=-44;bias1[192]=-117;bias1[193]=29;bias1[194]=-54;bias1[195]=-37;bias1[196]=-50;bias1[197]=12;bias1[198]=-27;bias1[199]=-63;


  end



endmodule
